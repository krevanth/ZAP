//////////////////////////////////////////////////////////////////////////////////
//                                                                              //                                    
//Copyright (C) 2016-2022 Revanth Kamaraj(krevanth) <revanth91kamaraj@gmail.com)//
//                                                                              // 
// This program is free software; you can redistribute it and/or                //
// modify it under the terms of the GNU General Public License                  //
// as published by the Free Software Foundation; either version 2               //
// of the License, or (at your option) any later version.                       //
//                                                                              //
// This program is distributed in the hope that it will be useful,              //
// but WITHOUT ANY WARRANTY; without even the implied warranty of               //
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the                //
// GNU General Public License for more details.                                 //
//                                                                              //
// You should have received a copy of the GNU General Public License            //
// along with this program; if not, write to the Free Software                  //
// Foundation, Inc., 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301,   //
// USA.                                                                         //
//                                                                              //
//////////////////////////////////////////////////////////////////////////////////
//                                                                              //
// Tag RAMs with single cycle clear. Finds the greatest use in TLBs.            //
//                                                                              //
//////////////////////////////////////////////////////////////////////////////////




module zap_mem_inv_block #(
        parameter DEPTH = 32,
        parameter WIDTH = 32   // Not including valid bit.
)(  


        input logic                           i_clk,
        input logic                           i_reset,
        input logic                           i_clken,

        // Write data.
        input logic   [WIDTH-1:0]             i_wdata,

        // Write and read enable.
        input logic                           i_wen, 

        // Invalidate entries in 1 cycle.
        input logic                           i_inv,

        // Read and write address.
        input logic   [$clog2(DEPTH)-1:0]     i_raddr, 
        input logic   [$clog2(DEPTH)-1:0]     i_waddr,

        // Read data and valid.
        output logic [WIDTH-1:0]              o_rdata,
        output logic                          o_rdav
);


logic [DEPTH-1:0]         dav_ff;
logic                     rdav;
logic                     rdav_st1;
logic [$clog2(DEPTH)-1:0] raddr_del;
logic                     sel_ff;

// Block RAM.
zap_ram_simple #(.WIDTH(WIDTH), .DEPTH(DEPTH)) u_ram_simple (
        .i_clk     ( i_clk ),
        .i_clken   ( i_clken ),

        .i_wr_en   ( i_wen ),

        .i_wr_data ( i_wdata ),
        .o_rd_data ( o_rdata ),

        .i_wr_addr ( i_waddr ),
        .i_rd_addr ( i_raddr )
);

// ----------------------------------------------------------------------------
// Stage 1
// ----------------------------------------------------------------------------

always_ff @ (posedge i_clk)
begin
        if ( i_reset | i_inv )
               dav_ff <= {DEPTH{1'd0}};
        else if ( i_wen && i_clken )
              dav_ff [ i_waddr ] <= 1'd1;
end

always @ ( posedge i_clk )
begin
        if ( i_reset || i_inv )
                rdav <= 1'd0;
        else if ( i_clken )
                rdav <= dav_ff [ i_raddr ];
end

always @ ( posedge i_clk )
begin
        if ( i_reset || i_inv )
                sel_ff <= 1'd0;
        else if ( i_clken )
                sel_ff <= i_raddr == i_waddr && i_wen;
end

always_ff @ ( posedge i_clk )
begin
        if ( i_reset || i_inv )
                raddr_del <= '0;
        else if ( i_clken )
                raddr_del <= i_raddr;
end

always_comb 
begin
        rdav_st1 = sel_ff ? 1'd1 : rdav;
end

// ----------------------------------------------------------------------------
// Stage 2
// ----------------------------------------------------------------------------

always_ff @ ( posedge i_clk )
begin
        if ( i_reset || i_inv )
                o_rdav <= 1'd0;
        else if  ( i_clken )
                o_rdav <= i_waddr == raddr_del && i_wen ? 1'd1 : rdav_st1;
end

endmodule // mem_inv_block.v

